`timescale 1ns / 1ps

module uart_rx(
    input clk50Mhz_i,
    input rst_i_n,
    input rx_i
    );
endmodule
