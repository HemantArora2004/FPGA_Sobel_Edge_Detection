`timescale 1ns / 1ps

module top_module(
    input clk,
    input uart_tx_out,
    output uart_rx_out,
    output led
    );
    
      
endmodule

   
